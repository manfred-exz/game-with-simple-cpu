module scinstmem_make_code_break_code (a,inst);   // instruction memory, rom
    input[31:0] a;                        // address
    output[31:0] inst;                    // instruction
    (* brom_map = "yes" *)
	reg[31:0] rom[0:124];

	assign inst = rom[a[8:2]];
    // rom[word_addr] = instruction
	assign rom[7'h0] = 32'h341d0ffc;
	assign rom[7'h1] = 32'h3c10a000;
	assign rom[7'h2] = 32'h3c11c000;
	assign rom[7'h3] = 32'h341200ff;
	assign rom[7'h4] = 32'h341300f0;
	assign rom[7'h5] = 32'h8e150000;
	assign rom[7'h6] = 32'h02a0402a;
	assign rom[7'h7] = 32'h1100fffd;
	assign rom[7'h8] = 32'h02b2b024;
	assign rom[7'h9] = 32'h340a00e0;
	assign rom[7'ha] = 32'h12cafffa;
	assign rom[7'hb] = 32'h12d3000d;
	assign rom[7'hc] = 32'h00162025;
	assign rom[7'hd] = 32'h34050001;
	assign rom[7'he] = 32'h0c000021;
	assign rom[7'hf] = 32'h1440fff5;
	assign rom[7'h10] = 32'h22d6fff2;
	assign rom[7'h11] = 32'h0016b080;
	assign rom[7'h12] = 32'h8ed40000;
	assign rom[7'h13] = 32'h36840000;
	assign rom[7'h14] = 32'h0c00004d;
	assign rom[7'h15] = 32'h34540000;
	assign rom[7'h16] = 32'hae340000;
	assign rom[7'h17] = 32'h22310004;
	assign rom[7'h18] = 32'h08000005;
	assign rom[7'h19] = 32'h8e150000;
	assign rom[7'h1a] = 32'h02a0402a;
	assign rom[7'h1b] = 32'h1100fffd;
	assign rom[7'h1c] = 32'h02b2b024;
	assign rom[7'h1d] = 32'h00162025;
	assign rom[7'h1e] = 32'h34050000;
	assign rom[7'h1f] = 32'h0c000021;
	assign rom[7'h20] = 32'h08000005;
	assign rom[7'h21] = 32'h34080058;
	assign rom[7'h22] = 32'h14880007;
	assign rom[7'h23] = 32'h14a00004;
	assign rom[7'h24] = 32'h3409014c;
	assign rom[7'h25] = 32'h8d2a0000;
	assign rom[7'h26] = 32'h394a0001;
	assign rom[7'h27] = 32'had2a0000;
	assign rom[7'h28] = 32'h34020001;
	assign rom[7'h29] = 32'h03e00008;
	assign rom[7'h2a] = 32'h34080012;
	assign rom[7'h2b] = 32'h10880003;
	assign rom[7'h2c] = 32'h34080059;
	assign rom[7'h2d] = 32'h10880001;
	assign rom[7'h2e] = 32'h08000033;
	assign rom[7'h2f] = 32'h34080144;
	assign rom[7'h30] = 32'had050000;
	assign rom[7'h31] = 32'h34020001;
	assign rom[7'h32] = 32'h03e00008;
	assign rom[7'h33] = 32'h34080014;
	assign rom[7'h34] = 32'h10880001;
	assign rom[7'h35] = 32'h0800003a;
	assign rom[7'h36] = 32'h34080140;
	assign rom[7'h37] = 32'had050000;
	assign rom[7'h38] = 32'h34020001;
	assign rom[7'h39] = 32'h03e00008;
	assign rom[7'h3a] = 32'h34080011;
	assign rom[7'h3b] = 32'h10880001;
	assign rom[7'h3c] = 32'h08000041;
	assign rom[7'h3d] = 32'h34080148;
	assign rom[7'h3e] = 32'had050000;
	assign rom[7'h3f] = 32'h34020001;
	assign rom[7'h40] = 32'h03e00008;
	assign rom[7'h41] = 32'h3408000e;
	assign rom[7'h42] = 32'h0088482a;
	assign rom[7'h43] = 32'h11200002;
	assign rom[7'h44] = 32'h34020001;
	assign rom[7'h45] = 32'h03e00008;
	assign rom[7'h46] = 32'h3408005d;
	assign rom[7'h47] = 32'h0104482a;
	assign rom[7'h48] = 32'h11200002;
	assign rom[7'h49] = 32'h34020001;
	assign rom[7'h4a] = 32'h03e00008;
	assign rom[7'h4b] = 32'h34020000;
	assign rom[7'h4c] = 32'h03e00008;
	assign rom[7'h4d] = 32'h34080026;
	assign rom[7'h4e] = 32'h34090061;
	assign rom[7'h4f] = 32'h0089502a;
	assign rom[7'h50] = 32'h0104582a;
	assign rom[7'h51] = 32'h11400029;
	assign rom[7'h52] = 32'h11600028;
	assign rom[7'h53] = 32'h23bdfff8;
	assign rom[7'h54] = 32'hafb20000;
	assign rom[7'h55] = 32'hafb30004;
	assign rom[7'h56] = 32'h3408014c;
	assign rom[7'h57] = 32'h8d120000;
	assign rom[7'h58] = 32'h34080144;
	assign rom[7'h59] = 32'h8d130000;
	assign rom[7'h5a] = 32'h3408003f;
	assign rom[7'h5b] = 32'h0088482a;
	assign rom[7'h5c] = 32'h1520000f;
	assign rom[7'h5d] = 32'h34080060;
	assign rom[7'h5e] = 32'h10880007;
	assign rom[7'h5f] = 32'h3408005b;
	assign rom[7'h60] = 32'h10880008;
	assign rom[7'h61] = 32'h3408005c;
	assign rom[7'h62] = 32'h10880006;
	assign rom[7'h63] = 32'h3408005d;
	assign rom[7'h64] = 32'h10880004;
	assign rom[7'h65] = 32'h08000072;
	assign rom[7'h66] = 32'h12600010;
	assign rom[7'h67] = 32'h2082001e;
	assign rom[7'h68] = 32'h08000078;
	assign rom[7'h69] = 32'h1260000d;
	assign rom[7'h6a] = 32'h20820020;
	assign rom[7'h6b] = 32'h08000078;
	assign rom[7'h6c] = 32'h1260000a;
	assign rom[7'h6d] = 32'h00044080;
	assign rom[7'h6e] = 32'h210800a4;
	assign rom[7'h6f] = 32'h8d090000;
	assign rom[7'h70] = 32'h35220000;
	assign rom[7'h71] = 32'h08000078;
	assign rom[7'h72] = 32'h02534026;
	assign rom[7'h73] = 32'h15000003;
	assign rom[7'h74] = 32'h34080020;
	assign rom[7'h75] = 32'h00881020;
	assign rom[7'h76] = 32'h08000078;
	assign rom[7'h77] = 32'h00801020;
	assign rom[7'h78] = 32'h8fb20000;
	assign rom[7'h79] = 32'h8fb30004;
	assign rom[7'h7a] = 32'h23bd0008;
	assign rom[7'h7b] = 32'h03e00008;
endmodule
