/************************************************
The Verilog HDL code example is from the book
Computer Principles and Design in Verilog HDL
by Yamin Li, published by A JOHN WILEY & SONS
************************************************/
module scinstmem_make_code_break_code (clk, a, inst); // instruction memory, rom
	input  clk;
	input  [31:0] a;                        	// address
	output reg [31:0] inst;                     	// instruction
//	wire   [31:0] rom [0:127];              	// rom cells: 64 words * 32 bits
	
	(* brom_map = "yes" *)
	reg [31:0] rom [0:127];
	
	always @(posedge clk)
		inst <= rom[a[8:2]];
	
//	assign inst = rom[a[8:2]];              	// use word address to read rom
	initial begin
		rom[7'd0] = 32'h341d0ffc;
		rom[7'd1] = 32'h3c10a000;
		rom[7'd2] = 32'h3c11c000;
		rom[7'd3] = 32'h341200ff;
		rom[7'd4] = 32'h341300f0;
		rom[7'd5] = 32'h8e150000;
		rom[7'd6] = 32'h02a0402a;
		rom[7'd7] = 32'h1100fffd;
		rom[7'd8] = 32'h02b2b024;
		rom[7'd9] = 32'h340a00e0;
		rom[7'd10] = 32'h12cafffa;
		rom[7'd11] = 32'h12d3000d;
		rom[7'd12] = 32'h00162025;
		rom[7'd13] = 32'h34050001;
		rom[7'd14] = 32'h0c000021;
		rom[7'd15] = 32'h1440fff5;
		rom[7'd16] = 32'h22d6fff2;
		rom[7'd17] = 32'h0016b080;
		rom[7'd18] = 32'h8ed40000;
		rom[7'd19] = 32'h36840000;
		rom[7'd20] = 32'h0c00004d;
		rom[7'd21] = 32'h34540000;
		rom[7'd22] = 32'hae340000;
		rom[7'd23] = 32'h22310004;
		rom[7'd24] = 32'h08000005;
		rom[7'd25] = 32'h8e150000;
		rom[7'd26] = 32'h02a0402a;
		rom[7'd27] = 32'h1100fffd;
		rom[7'd28] = 32'h02b2b024;
		rom[7'd29] = 32'h00162025;
		rom[7'd30] = 32'h34050000;
		rom[7'd31] = 32'h0c000021;
		rom[7'd32] = 32'h08000005;
		rom[7'd33] = 32'h34080058;
		rom[7'd34] = 32'h14880007;
		rom[7'd35] = 32'h14a00004;
		rom[7'd36] = 32'h3409014c;
		rom[7'd37] = 32'h8d2a0000;
		rom[7'd38] = 32'h394a0001;
		rom[7'd39] = 32'had2a0000;
		rom[7'd40] = 32'h34020001;
		rom[7'd41] = 32'h03e00008;
		rom[7'd42] = 32'h34080012;
		rom[7'd43] = 32'h10880003;
		rom[7'd44] = 32'h34080059;
		rom[7'd45] = 32'h10880001;
		rom[7'd46] = 32'h08000033;
		rom[7'd47] = 32'h34080144;
		rom[7'd48] = 32'had050000;
		rom[7'd49] = 32'h34020001;
		rom[7'd50] = 32'h03e00008;
		rom[7'd51] = 32'h34080014;
		rom[7'd52] = 32'h10880001;
		rom[7'd53] = 32'h0800003a;
		rom[7'd54] = 32'h34080140;
		rom[7'd55] = 32'had050000;
		rom[7'd56] = 32'h34020001;
		rom[7'd57] = 32'h03e00008;
		rom[7'd58] = 32'h34080011;
		rom[7'd59] = 32'h10880001;
		rom[7'd60] = 32'h08000041;
		rom[7'd61] = 32'h34080148;
		rom[7'd62] = 32'had050000;
		rom[7'd63] = 32'h34020001;
		rom[7'd64] = 32'h03e00008;
		rom[7'd65] = 32'h3408000e;
		rom[7'd66] = 32'h0088482a;
		rom[7'd67] = 32'h11200002;
		rom[7'd68] = 32'h34020001;
		rom[7'd69] = 32'h03e00008;
		rom[7'd70] = 32'h3408005d;
		rom[7'd71] = 32'h0104482a;
		rom[7'd72] = 32'h11200002;
		rom[7'd73] = 32'h34020001;
		rom[7'd74] = 32'h03e00008;
		rom[7'd75] = 32'h34020000;
		rom[7'd76] = 32'h03e00008;
		rom[7'd77] = 32'h34080026;
		rom[7'd78] = 32'h34090061;
		rom[7'd79] = 32'h0089502a;
		rom[7'd80] = 32'h0104582a;
		rom[7'd81] = 32'h11400029;
		rom[7'd82] = 32'h11600028;
		rom[7'd83] = 32'h23bdfff8;
		rom[7'd84] = 32'hafb20000;
		rom[7'd85] = 32'hafb30004;
		rom[7'd86] = 32'h3408014c;
		rom[7'd87] = 32'h8d120000;
		rom[7'd88] = 32'h34080144;
		rom[7'd89] = 32'h8d130000;
		rom[7'd90] = 32'h3408003f;
		rom[7'd91] = 32'h0088482a;
		rom[7'd92] = 32'h1520000f;
		rom[7'd93] = 32'h34080060;
		rom[7'd94] = 32'h10880007;
		rom[7'd95] = 32'h3408005b;
		rom[7'd96] = 32'h10880008;
		rom[7'd97] = 32'h3408005c;
		rom[7'd98] = 32'h10880006;
		rom[7'd99] = 32'h3408005d;
		rom[7'd100] = 32'h10880004;
		rom[7'd101] = 32'h08000072;
		rom[7'd102] = 32'h12600010;
		rom[7'd103] = 32'h2082001e;
		rom[7'd104] = 32'h08000078;
		rom[7'd105] = 32'h1260000d;
		rom[7'd106] = 32'h20820020;
		rom[7'd107] = 32'h08000078;
		rom[7'd108] = 32'h1260000a;
		rom[7'd109] = 32'h00044080;
		rom[7'd110] = 32'h210800a4;
		rom[7'd111] = 32'h8d090000;
		rom[7'd112] = 32'h35220000;
		rom[7'd113] = 32'h08000078;
		rom[7'd114] = 32'h02534026;
		rom[7'd115] = 32'h15000003;
		rom[7'd116] = 32'h34080020;
		rom[7'd117] = 32'h00881020;
		rom[7'd118] = 32'h08000078;
		rom[7'd119] = 32'h00801020;
		rom[7'd120] = 32'h8fb20000;
		rom[7'd121] = 32'h8fb30004;
		rom[7'd122] = 32'h23bd0008;
		rom[7'd123] = 32'h03e00008;
	end


//rom[7'd0] = 32'h341d0ffc;
//rom[7'd1] = 32'h3c10a000;
//rom[7'd2] = 32'h3c11c000;
//rom[7'd3] = 32'h341200ff;
//rom[7'd4] = 32'h341300f0;
//rom[7'd5] = 32'h34170001;
//rom[7'd6] = 32'h8e150000;
//rom[7'd7] = 32'h02a0402a;
//rom[7'd8] = 32'h1100fffd;
//rom[7'd9] = 32'h02b2b024;
//rom[7'd10] = 32'h340a00e0;
//rom[7'd11] = 32'h12cafffa;
//rom[7'd12] = 32'h00162025;
//rom[7'd13] = 32'h34050001;
//rom[7'd14] = 32'h0c000022;
//rom[7'd15] = 32'h1440fff6;
//rom[7'd16] = 32'h12d30009;
//rom[7'd17] = 32'h22d6fff2;
//rom[7'd18] = 32'h0016b080;
//rom[7'd19] = 32'h8ed40000;
//rom[7'd20] = 32'h36840000;
//rom[7'd21] = 32'h0c000041;
//rom[7'd22] = 32'h34540000;
//rom[7'd23] = 32'hae340000;
//rom[7'd24] = 32'h22310004;
//rom[7'd25] = 32'h08000006;
//rom[7'd26] = 32'h8e150000;
//rom[7'd27] = 32'h02a0402a;
//rom[7'd28] = 32'h1100fffd;
//rom[7'd29] = 32'h02b2b024;
//rom[7'd30] = 32'h00162025;
//rom[7'd31] = 32'h34050000;
//rom[7'd32] = 32'h0c000022;
//rom[7'd33] = 32'h08000006;
//rom[7'd34] = 32'h34080058;
//rom[7'd35] = 32'h14880004;
//rom[7'd36] = 32'h3409014c;
//rom[7'd37] = 32'h8d2a0000;
//rom[7'd38] = 32'h394a0001;
//rom[7'd39] = 32'had2a0000;
//rom[7'd40] = 32'h34080012;
//rom[7'd41] = 32'h10880003;
//rom[7'd42] = 32'h34080059;
//rom[7'd43] = 32'h10880001;
//rom[7'd44] = 32'h08000031;
//rom[7'd45] = 32'h34080144;
//rom[7'd46] = 32'had050000;
//rom[7'd47] = 32'h34020001;
//rom[7'd48] = 32'h03e00008;
//rom[7'd49] = 32'h34080014;
//rom[7'd50] = 32'h10880001;
//rom[7'd51] = 32'h08000038;
//rom[7'd52] = 32'h34080140;
//rom[7'd53] = 32'had050000;
//rom[7'd54] = 32'h34020001;
//rom[7'd55] = 32'h03e00008;
//rom[7'd56] = 32'h34080011;
//rom[7'd57] = 32'h10880001;
//rom[7'd58] = 32'h0800003f;
//rom[7'd59] = 32'h34080148;
//rom[7'd60] = 32'had050000;
//rom[7'd61] = 32'h34020001;
//rom[7'd62] = 32'h03e00008;
//rom[7'd63] = 32'h34020000;
//rom[7'd64] = 32'h03e00008;
//rom[7'd65] = 32'h34080026;
//rom[7'd66] = 32'h34090061;
//rom[7'd67] = 32'h0089502a;
//rom[7'd68] = 32'h0104582a;
//rom[7'd69] = 32'h11400023;
//rom[7'd70] = 32'h11600022;
//rom[7'd71] = 32'h23bdfff8;
//rom[7'd72] = 32'hafb20000;
//rom[7'd73] = 32'hafb30004;
//rom[7'd74] = 32'h3408014c;
//rom[7'd75] = 32'h8d120000;
//rom[7'd76] = 32'h34080144;
//rom[7'd77] = 32'h8d130000;
//rom[7'd78] = 32'h3408003f;
//rom[7'd79] = 32'h0088482a;
//rom[7'd80] = 32'h15200009;
//rom[7'd81] = 32'h3508005a;
//rom[7'd82] = 32'h0104482a;
//rom[7'd83] = 32'h15200006;
//rom[7'd84] = 32'h01004020;
//rom[7'd85] = 32'h01004020;
//rom[7'd86] = 32'h01004020;
//rom[7'd87] = 32'h01004020;
//rom[7'd88] = 32'h01004020;
//rom[7'd89] = 32'h08000060;
//rom[7'd90] = 32'h1260000a;
//rom[7'd91] = 32'h00044080;
//rom[7'd92] = 32'h210800a4;
//rom[7'd93] = 32'h8d090000;
//rom[7'd94] = 32'h35220000;
//rom[7'd95] = 32'h08000066;
//rom[7'd96] = 32'h02534026;
//rom[7'd97] = 32'h15000003;
//rom[7'd98] = 32'h34080020;
//rom[7'd99] = 32'h00881020;
//rom[7'd100] = 32'h08000066;
//rom[7'd101] = 32'h00801020;
//rom[7'd102] = 32'h8fb20000;
//rom[7'd103] = 32'h8fb30004;
//rom[7'd104] = 32'h23bd0008;
//rom[7'd105] = 32'h03e00008;

	
//	 rom[word_addr] = instruction
//	assign rom[7'd0] = 32'h341d0400;
//	assign rom[7'd1] = 32'h3c10a000;
//	assign rom[7'd2] = 32'h3c11c000;
//	assign rom[7'd3] = 32'h341200ff;
//	assign rom[7'd4] = 32'h341300f0;
//	assign rom[7'd5] = 32'h34170001;
//	assign rom[7'd6] = 32'h8e150000;
//	assign rom[7'd7] = 32'h02a0402a;
//	assign rom[7'd8] = 32'h1100fffd;
//	assign rom[7'd9] = 32'h02b2b024;
//	assign rom[7'd10] = 32'h340a00e0;
//	assign rom[7'd11] = 32'h12cafffa;
//	assign rom[7'd12] = 32'h00162025;
//	assign rom[7'd13] = 32'h34050001;
//	assign rom[7'd14] = 32'h0c000022;
//	assign rom[7'd15] = 32'h1440fff6;
//	assign rom[7'd16] = 32'h12d30009;
//	assign rom[7'd17] = 32'h22d6fff2;
//	assign rom[7'd18] = 32'h0016b080;
//	assign rom[7'd19] = 32'h8ed40000;
//	assign rom[7'd20] = 32'h36840000;
//	assign rom[7'd21] = 32'h0c000041;
//	assign rom[7'd22] = 32'h34540000;
//	assign rom[7'd23] = 32'hae340000;
//	assign rom[7'd24] = 32'h22310004;
//	assign rom[7'd25] = 32'h08000006;
//	assign rom[7'd26] = 32'h8e150000;
//	assign rom[7'd27] = 32'h02a0402a;
//	assign rom[7'd28] = 32'h1100fffd;
//	assign rom[7'd29] = 32'h02b2b024;
//	assign rom[7'd30] = 32'h00162025;
//	assign rom[7'd31] = 32'h34050000;
//	assign rom[7'd32] = 32'h0c000022;
//	assign rom[7'd33] = 32'h08000006;
//	assign rom[7'd34] = 32'h34080058;
//	assign rom[7'd35] = 32'h14880004;
//	assign rom[7'd36] = 32'h3409014c;
//	assign rom[7'd37] = 32'h8d2a0000;
//	assign rom[7'd38] = 32'h394a0001;
//	assign rom[7'd39] = 32'had2a0000;
//	assign rom[7'd40] = 32'h34080012;
//	assign rom[7'd41] = 32'h10880003;
//	assign rom[7'd42] = 32'h34080059;
//	assign rom[7'd43] = 32'h10880001;
//	assign rom[7'd44] = 32'h08000031;
//	assign rom[7'd45] = 32'h34080144;
//	assign rom[7'd46] = 32'had050000;
//	assign rom[7'd47] = 32'h34020001;
//	assign rom[7'd48] = 32'h03e00008;
//	assign rom[7'd49] = 32'h34080014;
//	assign rom[7'd50] = 32'h10880001;
//	assign rom[7'd51] = 32'h08000038;
//	assign rom[7'd52] = 32'h34080140;
//	assign rom[7'd53] = 32'had050000;
//	assign rom[7'd54] = 32'h34020001;
//	assign rom[7'd55] = 32'h03e00008;
//	assign rom[7'd56] = 32'h34080011;
//	assign rom[7'd57] = 32'h10880001;
//	assign rom[7'd58] = 32'h0800003f;
//	assign rom[7'd59] = 32'h34080148;
//	assign rom[7'd60] = 32'had050000;
//	assign rom[7'd61] = 32'h34020001;
//	assign rom[7'd62] = 32'h03e00008;
//	assign rom[7'd63] = 32'h34020000;
//	assign rom[7'd64] = 32'h03e00008;
//	assign rom[7'd65] = 32'h34080026;
//	assign rom[7'd66] = 32'h34090061;
//	assign rom[7'd67] = 32'h0089502a;
//	assign rom[7'd68] = 32'h0104582a;
//	assign rom[7'd69] = 32'h1140001c;
//	assign rom[7'd70] = 32'h1160001b;
//	assign rom[7'd71] = 32'h23bdfff8;
//	assign rom[7'd72] = 32'hafb00000;
//	assign rom[7'd73] = 32'hafb10004;
//	assign rom[7'd74] = 32'h3408014c;
//	assign rom[7'd75] = 32'h8d100000;
//	assign rom[7'd76] = 32'h34080144;
//	assign rom[7'd77] = 32'h8d110000;
//	assign rom[7'd78] = 32'h3508003f;
//	assign rom[7'd79] = 32'h0088482a;
//	assign rom[7'd80] = 32'h15200004;
//	assign rom[7'd81] = 32'h3508005a;
//	assign rom[7'd82] = 32'h0104482a;
//	assign rom[7'd83] = 32'h15200001;
//	assign rom[7'd84] = 32'h0800005b;
//	assign rom[7'd85] = 32'h12200008;
//	assign rom[7'd86] = 32'h00044080;
//	assign rom[7'd87] = 32'h210800a4;
//	assign rom[7'd88] = 32'h8d090000;
//	assign rom[7'd89] = 32'h35220000;
//	assign rom[7'd90] = 32'h0800005f;
//	assign rom[7'd91] = 32'h02114026;
//	assign rom[7'd92] = 32'h15000001;
//	assign rom[7'd93] = 32'h20820020;
//	assign rom[7'd94] = 32'h00801020;
//	assign rom[7'd95] = 32'h8fb00000;
//	assign rom[7'd96] = 32'h8fb10004;
//	assign rom[7'd97] = 32'h23bd0008;
//	assign rom[7'd98] = 32'h03e00008;

//
//	assign rom[6'd0] = 32'h341d0200;
//	assign rom[6'd1] = 32'h3c10a000;
//	assign rom[6'd2] = 32'h3c11c000;
//	assign rom[6'd3] = 32'h341200ff;
//	assign rom[6'd4] = 32'h341300f0;
//	assign rom[6'd5] = 32'h34170001;
//	assign rom[6'd6] = 32'h8e150000;
//	assign rom[6'd7] = 32'h02a0402a;
//	assign rom[6'd8] = 32'h1100fffd;
//	assign rom[6'd9] = 32'h02b2b024;
//	assign rom[6'd10] = 32'h340a00e0;
//	assign rom[6'd11] = 32'h12cafffa;
//	assign rom[6'd12] = 32'h00162025;
//	assign rom[6'd13] = 32'h34050001;
//	assign rom[6'd14] = 32'h0c00001f;
//	assign rom[6'd15] = 32'h1440fff6;
//	assign rom[6'd16] = 32'h12d30006;
//	assign rom[6'd17] = 32'h22d6fff2;
//	assign rom[6'd18] = 32'h0016b080;
//	assign rom[6'd19] = 32'h8ed40000;
//	assign rom[6'd20] = 32'hae340000;
//	assign rom[6'd21] = 32'h22310004;
//	assign rom[6'd22] = 32'h08000006;
//	assign rom[6'd23] = 32'h8e150000;
//	assign rom[6'd24] = 32'h02a0402a;
//	assign rom[6'd25] = 32'h1100fffd;
//	assign rom[6'd26] = 32'h02b2b024;
//	assign rom[6'd27] = 32'h00162025;
//	assign rom[6'd28] = 32'h34050000;
//	assign rom[6'd29] = 32'h0c00001f;
//	assign rom[6'd30] = 32'h08000006;
//	assign rom[6'd31] = 32'h34080012;
//	assign rom[6'd32] = 32'h10880003;
//	assign rom[6'd33] = 32'h34080059;
//	assign rom[6'd34] = 32'h10880001;
//	assign rom[6'd35] = 32'h08000028;
//	assign rom[6'd36] = 32'h34080144;
//	assign rom[6'd37] = 32'had050000;
//	assign rom[6'd38] = 32'h34020001;
//	assign rom[6'd39] = 32'h03e00008;
//	assign rom[6'd40] = 32'h34080014;
//	assign rom[6'd41] = 32'h10880001;
//	assign rom[6'd42] = 32'h0800002f;
//	assign rom[6'd43] = 32'h34080140;
//	assign rom[6'd44] = 32'had050000;
//	assign rom[6'd45] = 32'h34020001;
//	assign rom[6'd46] = 32'h03e00008;
//	assign rom[6'd47] = 32'h34080011;
//	assign rom[6'd48] = 32'h10880001;
//	assign rom[6'd49] = 32'h08000036;
//	assign rom[6'd50] = 32'h34080148;
//	assign rom[6'd51] = 32'had050000;
//	assign rom[6'd52] = 32'h34020001;
//	assign rom[6'd53] = 32'h03e00008;
//	assign rom[6'd54] = 32'h34020000;
//	assign rom[6'd55] = 32'h03e00008;


//	assign rom[6'h00] = 32'b00111100000000111100000000000000;
//	assign rom[6'h01] = 32'b00111100000001001010000000000000;
//	assign rom[6'h02] = 32'b10001100100001010000000000000000;
//	assign rom[6'h03] = 32'b00110000101001100000000100000000;
//	assign rom[6'h04] = 32'b00010000110000001111111111111101;
//	assign rom[6'h05] = 32'b00110000101001100000000011111111;
//	assign rom[6'h06] = 32'b00000000000001100010100100000010;
//	assign rom[6'h07] = 32'b00100000101001111111111111110110;
//	assign rom[6'h08] = 32'b00000000000001110011111111000010;
//	assign rom[6'h09] = 32'b00010000111000000000000000000010;
//	assign rom[6'h0a] = 32'b00100000101001010000000000110000;
//	assign rom[6'h0b] = 32'b00001000000000000000000000001101;
//	assign rom[6'h0c] = 32'b00100000101001010000000000110111;
//	assign rom[6'h0d] = 32'b00001100000000000000000000011001;
//	assign rom[6'h0e] = 32'b00110000110001010000000000001111;
//	assign rom[6'h0f] = 32'b00100000101001111111111111110110;
//	assign rom[6'h10] = 32'b00000000000001110011111111000010;
//	assign rom[6'h11] = 32'b00010000111000000000000000000010;
//	assign rom[6'h12] = 32'b00100000101001010000000000110000;
//	assign rom[6'h13] = 32'b00001000000000000000000000010101;
//	assign rom[6'h14] = 32'b00100000101001010000000000110111;
//	assign rom[6'h15] = 32'b00001100000000000000000000011001;
//	assign rom[6'h16] = 32'b00100000000001010000000000100000;
//	assign rom[6'h17] = 32'b00001100000000000000000000011001;
//	assign rom[6'h18] = 32'b00001000000000000000000000000010;
//	assign rom[6'h19] = 32'b10101100011001010000000000000000;
//	assign rom[6'h1a] = 32'b00100000011000110000000000000100;
//	assign rom[6'h1b] = 32'b00000011111000000000000000001000;
//	assign rom[6'h1c] = 32'b00000000000000000000000000000000;
//	assign rom[6'h1d] = 32'b00000000000000000000000000000000;
//	assign rom[6'h1e] = 32'b00000000000000000000000000000000;
//	assign rom[6'h1f] = 32'b00000000000000000000000000000000;
endmodule
