module scinstmem_make_code_break_code (a,inst);	// instruction memory, rom
	input	[31:0]  a;								// address
	output	[31:0] inst;						// instruction

	(* brom_map = "yes" *)
	reg[31:0] rom[0:257];

	assign inst = rom[a[10:2]];

	initial begin
		rom[9'h0] = 32'h241d0ffc;
		rom[9'h1] = 32'h8c0801b0;
		rom[9'h2] = 32'h0800004d;
		rom[9'h3] = 32'h8c1801ac;
		rom[9'h4] = 32'h83020000;
		rom[9'h5] = 32'h23180001;
		rom[9'h6] = 32'hac1801ac;
		rom[9'h7] = 32'h03e00008;
		rom[9'h8] = 32'h23bdfff8;
		rom[9'h9] = 32'hafb00000;
		rom[9'ha] = 32'hafbf0004;
		rom[9'hb] = 32'h00048021;
		rom[9'hc] = 32'h8c0401a4;
		rom[9'hd] = 32'h8c0501a8;
		rom[9'he] = 32'h0c000016;
		rom[9'hf] = 32'h00000000;
		rom[9'h10] = 32'hac500000;
		rom[9'h11] = 32'h00000000;
		rom[9'h12] = 32'h8fbf0004;
		rom[9'h13] = 32'h8fb00000;
		rom[9'h14] = 32'h23bd0008;
		rom[9'h15] = 32'h03e00008;
		rom[9'h16] = 32'h3c01c000;
		rom[9'h17] = 32'h34220000;
		rom[9'h18] = 32'h00054200;
		rom[9'h19] = 32'h00054980;
		rom[9'h1a] = 32'h00481020;
		rom[9'h1b] = 32'h00491020;
		rom[9'h1c] = 32'h00045080;
		rom[9'h1d] = 32'h004a1020;
		rom[9'h1e] = 32'h03e00008;
		rom[9'h1f] = 32'h8c0801a8;
		rom[9'h20] = 32'h2409003b;
		rom[9'h21] = 32'h15090004;
		rom[9'h22] = 32'h24080000;
		rom[9'h23] = 32'hac0801a8;
		rom[9'h24] = 32'h00081021;
		rom[9'h25] = 32'h03e00008;
		rom[9'h26] = 32'h21080001;
		rom[9'h27] = 32'hac0801a8;
		rom[9'h28] = 32'h00081021;
		rom[9'h29] = 32'h03e00008;
		rom[9'h2a] = 32'h23bdfffc;
		rom[9'h2b] = 32'hafbf0000;
		rom[9'h2c] = 32'h0c000035;
		rom[9'h2d] = 32'h2409004f;
		rom[9'h2e] = 32'h0122402a;
		rom[9'h2f] = 32'h11000001;
		rom[9'h30] = 32'h2042ffb1;
		rom[9'h31] = 32'hac0201a4;
		rom[9'h32] = 32'h8fbf0000;
		rom[9'h33] = 32'h23bd0004;
		rom[9'h34] = 32'h03e00008;
		rom[9'h35] = 32'h3c011000;
		rom[9'h36] = 32'h34380100;
		rom[9'h37] = 32'h8f020000;
		rom[9'h38] = 32'h2408007f;
		rom[9'h39] = 32'h00481024;
		rom[9'h3a] = 32'h03e00008;
		rom[9'h3b] = 32'h23bdfff4;
		rom[9'h3c] = 32'hafb10008;
		rom[9'h3d] = 32'hafbf0004;
		rom[9'h3e] = 32'hafb00000;
		rom[9'h3f] = 32'h00042821;
		rom[9'h40] = 32'h24100000;
		rom[9'h41] = 32'h24110050;
		rom[9'h42] = 32'h00102021;
		rom[9'h43] = 32'h0c000016;
		rom[9'h44] = 32'hac400000;
		rom[9'h45] = 32'h12110002;
		rom[9'h46] = 32'h22100001;
		rom[9'h47] = 32'h08000042;
		rom[9'h48] = 32'h8fb10008;
		rom[9'h49] = 32'h8fb00000;
		rom[9'h4a] = 32'h8fbf0004;
		rom[9'h4b] = 32'h23bd0008;
		rom[9'h4c] = 32'h03e00008;
		rom[9'h4d] = 32'h24020000;
		rom[9'h4e] = 32'h0c000083;
		rom[9'h4f] = 32'h8c1801b4;
		rom[9'h50] = 32'h83080000;
		rom[9'h51] = 32'h15000003;
		rom[9'h52] = 32'h23180001;
		rom[9'h53] = 32'hac1801b4;
		rom[9'h54] = 32'h0800004f;
		rom[9'h55] = 32'h11020001;
		rom[9'h56] = 32'h08000066;
		rom[9'h57] = 32'h8c0901ac;
		rom[9'h58] = 32'h8c0a01b4;
		rom[9'h59] = 32'h112a000c;
		rom[9'h5a] = 32'h21480001;
		rom[9'h5b] = 32'hac0801b4;
		rom[9'h5c] = 32'h8c0401b8;
		rom[9'h5d] = 32'h0c00003b;
		rom[9'h5e] = 32'h8c0801b8;
		rom[9'h5f] = 32'h2409003b;
		rom[9'h60] = 32'h11090001;
		rom[9'h61] = 32'h08000064;
		rom[9'h62] = 32'hac0001b8;
		rom[9'h63] = 32'h08000066;
		rom[9'h64] = 32'h21080001;
		rom[9'h65] = 32'hac0801b8;
		rom[9'h66] = 32'h3c010100;
		rom[9'h67] = 32'h34290000;
		rom[9'h68] = 32'h3c011000;
		rom[9'h69] = 32'h34380100;
		rom[9'h6a] = 32'h8c0801a0;
		rom[9'h6b] = 32'h01094024;
		rom[9'h6c] = 32'h11000003;
		rom[9'h6d] = 32'h8f0a0000;
		rom[9'h6e] = 32'hac0a01a0;
		rom[9'h6f] = 32'h0800004d;
		rom[9'h70] = 32'h8f080000;
		rom[9'h71] = 32'hac0801a0;
		rom[9'h72] = 32'h01094024;
		rom[9'h73] = 32'h1100ffd9;
		rom[9'h74] = 32'h08000075;
		rom[9'h75] = 32'h0c000003;
		rom[9'h76] = 32'h00024021;
		rom[9'h77] = 32'h24090003;
		rom[9'h78] = 32'h11280009;
		rom[9'h79] = 32'h15000002;
		rom[9'h7a] = 32'h0c00002a;
		rom[9'h7b] = 32'h08000075;
		rom[9'h7c] = 32'h00082021;
		rom[9'h7d] = 32'h0c000008;
		rom[9'h7e] = 32'h0c00001f;
		rom[9'h7f] = 32'h00022021;
		rom[9'h80] = 32'h0c00003b;
		rom[9'h81] = 32'h0800004d;
		rom[9'h82] = 32'h08000082;
		rom[9'h83] = 32'h23bdfffc;
		rom[9'h84] = 32'hafbf0000;
		rom[9'h85] = 32'h3c10a000;
		rom[9'h86] = 32'h3c11c000;
		rom[9'h87] = 32'h341200ff;
		rom[9'h88] = 32'h341300f0;
		rom[9'h89] = 32'h8e150000;
		rom[9'h8a] = 32'h02a0402a;
		rom[9'h8b] = 32'h11000017;
		rom[9'h8c] = 32'h02b2b024;
		rom[9'h8d] = 32'h340a00e0;
		rom[9'h8e] = 32'h12cafff4;
		rom[9'h8f] = 32'h12d3000c;
		rom[9'h90] = 32'h00162025;
		rom[9'h91] = 32'h34050001;
		rom[9'h92] = 32'h0c0000a6;
		rom[9'h93] = 32'h1440000f;
		rom[9'h94] = 32'h22d6fff2;
		rom[9'h95] = 32'h0016b080;
		rom[9'h96] = 32'h8ed40000;
		rom[9'h97] = 32'h36840000;
		rom[9'h98] = 32'h0c0000d2;
		rom[9'h99] = 32'h34540000;
		rom[9'h9a] = 32'h00141021;
		rom[9'h9b] = 32'h080000a3;
		rom[9'h9c] = 32'h8e150000;
		rom[9'h9d] = 32'h02a0402a;
		rom[9'h9e] = 32'h1100fffd;
		rom[9'h9f] = 32'h02b2b024;
		rom[9'ha0] = 32'h00162025;
		rom[9'ha1] = 32'h34050000;
		rom[9'ha2] = 32'h0c0000a6;
		rom[9'ha3] = 32'h8fbf0000;
		rom[9'ha4] = 32'h23bd0004;
		rom[9'ha5] = 32'h03e00008;
		rom[9'ha6] = 32'h34080058;
		rom[9'ha7] = 32'h14880007;
		rom[9'ha8] = 32'h14a00004;
		rom[9'ha9] = 32'h340901c8;
		rom[9'haa] = 32'h8d2a0000;
		rom[9'hab] = 32'h394a0001;
		rom[9'hac] = 32'had2a0000;
		rom[9'had] = 32'h34020001;
		rom[9'hae] = 32'h03e00008;
		rom[9'haf] = 32'h34080012;
		rom[9'hb0] = 32'h10880003;
		rom[9'hb1] = 32'h34080059;
		rom[9'hb2] = 32'h10880001;
		rom[9'hb3] = 32'h080000b8;
		rom[9'hb4] = 32'h340801c0;
		rom[9'hb5] = 32'had050000;
		rom[9'hb6] = 32'h34020001;
		rom[9'hb7] = 32'h03e00008;
		rom[9'hb8] = 32'h34080014;
		rom[9'hb9] = 32'h10880001;
		rom[9'hba] = 32'h080000bf;
		rom[9'hbb] = 32'h340801bc;
		rom[9'hbc] = 32'had050000;
		rom[9'hbd] = 32'h34020001;
		rom[9'hbe] = 32'h03e00008;
		rom[9'hbf] = 32'h34080011;
		rom[9'hc0] = 32'h10880001;
		rom[9'hc1] = 32'h080000c6;
		rom[9'hc2] = 32'h340801c4;
		rom[9'hc3] = 32'had050000;
		rom[9'hc4] = 32'h34020001;
		rom[9'hc5] = 32'h03e00008;
		rom[9'hc6] = 32'h3408000e;
		rom[9'hc7] = 32'h0088482a;
		rom[9'hc8] = 32'h11200002;
		rom[9'hc9] = 32'h34020001;
		rom[9'hca] = 32'h03e00008;
		rom[9'hcb] = 32'h3408005d;
		rom[9'hcc] = 32'h0104482a;
		rom[9'hcd] = 32'h11200002;
		rom[9'hce] = 32'h34020001;
		rom[9'hcf] = 32'h03e00008;
		rom[9'hd0] = 32'h34020000;
		rom[9'hd1] = 32'h03e00008;
		rom[9'hd2] = 32'h34080026;
		rom[9'hd3] = 32'h34090061;
		rom[9'hd4] = 32'h0089502a;
		rom[9'hd5] = 32'h0104582a;
		rom[9'hd6] = 32'h11400029;
		rom[9'hd7] = 32'h11600028;
		rom[9'hd8] = 32'h23bdfff8;
		rom[9'hd9] = 32'hafb20000;
		rom[9'hda] = 32'hafb30004;
		rom[9'hdb] = 32'h340801c8;
		rom[9'hdc] = 32'h8d120000;
		rom[9'hdd] = 32'h340801c0;
		rom[9'hde] = 32'h8d130000;
		rom[9'hdf] = 32'h3408003f;
		rom[9'he0] = 32'h0088482a;
		rom[9'he1] = 32'h1520000f;
		rom[9'he2] = 32'h34080060;
		rom[9'he3] = 32'h10880007;
		rom[9'he4] = 32'h3408005b;
		rom[9'he5] = 32'h10880008;
		rom[9'he6] = 32'h3408005c;
		rom[9'he7] = 32'h10880006;
		rom[9'he8] = 32'h3408005d;
		rom[9'he9] = 32'h10880004;
		rom[9'hea] = 32'h080000f7;
		rom[9'heb] = 32'h12600010;
		rom[9'hec] = 32'h2082001e;
		rom[9'hed] = 32'h080000fd;
		rom[9'hee] = 32'h1260000d;
		rom[9'hef] = 32'h20820020;
		rom[9'hf0] = 32'h080000fd;
		rom[9'hf1] = 32'h1260000a;
		rom[9'hf2] = 32'h00044080;
		rom[9'hf3] = 32'h210800a4;
		rom[9'hf4] = 32'h8d090000;
		rom[9'hf5] = 32'h35220000;
		rom[9'hf6] = 32'h080000fd;
		rom[9'hf7] = 32'h02534026;
		rom[9'hf8] = 32'h15000003;
		rom[9'hf9] = 32'h34080020;
		rom[9'hfa] = 32'h00881020;
		rom[9'hfb] = 32'h080000fd;
		rom[9'hfc] = 32'h00801020;
		rom[9'hfd] = 32'h8fb20000;
		rom[9'hfe] = 32'h8fb30004;
		rom[9'hff] = 32'h23bd0008;
		rom[9'h100] = 32'h03e00008;
	end

endmodule
