/************************************************
  The Verilog HDL code example is from the book
  Computer Principles and Design in Verilog HDL
  by Yamin Li, published by A JOHN WILEY & SONS
************************************************/
module single_cycle_cpu_io (clk,clrn,pc,inst,m_addr,m_write,m_read,d_f_mem,d_t_mem
                            ); 								// cpu kbd i/o
	input  clk, clrn;                                   	// clock and reset
	//[inst] read from mem
	input  [31:0] 	inst;                                 	// instruction
	//[data address/enable] for mem space
	output [31:0] 	m_addr;                               	// mem or i/o addr
	output 			m_write;
	output 			m_read;
	//[data] from/to mem
	input  [31:0] 	d_f_mem;                              	// load data
	output [31:0] 	d_t_mem;                              	// store data
	
	output [31:0] 	pc;                                   	// program counter
	
	
	// control signals
	reg           wreg = 0;                                 // write regfile
	reg           wmem = 0,rmem = 0;                        // write/read memory
	reg    [31:0] alu_out = 0;                              // alu output
	reg     [4:0] dest_rn = 0;                              // dest reg number
	reg    [31:0] next_pc = 0;                              // next pc
	wire   [31:0] pc_plus_4 = pc + 4;                   	// pc + 4
	
	// instruction format
	wire  [05:00] opcode = inst[31:26];
	wire  [04:00] rs     = inst[25:21];
	wire  [04:00] rt     = inst[20:16];
	wire  [04:00] rd     = inst[15:11];
	wire  [04:00] sa     = inst[10:06];
	wire  [05:00] func   = inst[05:00];
	wire  [15:00] imm    = inst[15:00];
	wire  [25:00] addr   = inst[25:00];
	wire          sign   = inst[15];
	wire  [31:00] offset = {{14{sign}},imm,2'b00};
	wire  [31:00] j_addr = {pc_plus_4[31:28],addr,2'b00};
	
	// instruction decode
	wire i_add  = (opcode == 6'h00) & (func == 6'h20);  // add
	wire i_sub  = (opcode == 6'h00) & (func == 6'h22);  // sub
	wire i_and  = (opcode == 6'h00) & (func == 6'h24);  // and
	wire i_or   = (opcode == 6'h00) & (func == 6'h25);  // or
	wire i_xor  = (opcode == 6'h00) & (func == 6'h26);  // xor
	wire i_sll  = (opcode == 6'h00) & (func == 6'h00);  // sll
	wire i_srl  = (opcode == 6'h00) & (func == 6'h02);  // srl
	wire i_sra  = (opcode == 6'h00) & (func == 6'h03);  // sra
	wire i_jr   = (opcode == 6'h00) & (func == 6'h08);  // jr
	wire i_addi = (opcode == 6'h08);                    // addi
	wire i_andi = (opcode == 6'h0c);                    // andi
	wire i_ori  = (opcode == 6'h0d);                    // ori
	wire i_xori = (opcode == 6'h0e);                    // xori
	wire i_lw   = (opcode == 6'h23);                    // lw
	wire i_sw   = (opcode == 6'h2b);                    // sw
	wire i_beq  = (opcode == 6'h04);                    // beq
	wire i_bne  = (opcode == 6'h05);                    // bne
	wire i_lui  = (opcode == 6'h0f);                    // lui
	wire i_j    = (opcode == 6'h02);                    // j
	wire i_jal  = (opcode == 6'h03);                    // jal
	
	wire i_slt  = (opcode == 6'h00) & (func == 6'h2a);	//slt
	wire i_slti = (opcode == 6'h0a);					//slti
	wire i_addiu= (opcode == 6'h09);
	wire i_addu = (opcode == 6'h00) & (func == 6'h21);	//addu
	
	wire i_lx = i_lb|i_lbu|i_lw;
	wire i_lb	= (opcode == 6'h20);					//lb
	wire i_lbu	= (opcode == 6'h24);					//lbu
	// sb: TO DO
//	wire i_sb	= (opcode == 6'h28);					//sb
	
//	wire signed [31:0]signed_a = a, signed_b = b;
	
	// pc
	reg [31:0] pc = -4;
	always @ (posedge clk or negedge clrn) begin
		if (!clrn) pc <= 0;
		else         pc <= next_pc;
	end
	
	
	// byte data or half-word data written to register file
//	wire [7:0]b_d_f_mem = d_f_mem[ m_addr[1:0] << 3 : m_addr[1:0] << 3 + 7];
	wire [7:0]b_d_f_mem = 	m_addr[1:0] == 2'b00 ? d_f_mem[7:0] : (
							m_addr[1:0] == 2'b01 ? d_f_mem[15:8]: (
							m_addr[1:0] == 2'b10 ? d_f_mem[23:16]: 
											   d_f_mem[31:24]
											   )
											   );
	
	// data written to register file
//	wire   [31:0] data_2_rf = i_lw ? d_f_mem : alu_out;
	wire   [31:0] data_2_rf = i_lb ? { {24{b_d_f_mem[7]}}, b_d_f_mem } : 
										(i_lbu ? {24'h0, b_d_f_mem} : 
											(i_lw ? d_f_mem : alu_out
											)
										);
	
	// register file
	reg    [31:0] regfile [1:31];                       // $1 - $31
	wire   [31:0] a = (rs==0) ? 0 : regfile[rs];        // read port
	wire   [31:0] b = (rt==0) ? 0 : regfile[rt];        // read port
	integer i;
	initial begin 
		for(i = 1; i < 32; i = i+1)
			regfile[i] = 32'h0;
	end
	
	always @ (posedge clk) begin
	  if (wreg && (dest_rn != 0)) begin
			regfile[dest_rn] <= data_2_rf;              // write port
	  end
	end
	
	// output signals
	assign m_read 	= rmem;
	assign m_write = wmem;
	assign d_t_mem =   b;                               // data to store
	// store byte: TO DO
//	assign d_t_mem =   i_sb ? 							
	assign m_addr  =   (i_lw|i_sw|i_lx) ? alu_out : 32'h0;                         // memory address
	

	// control signals, will be combinational circuit
	always @(*) begin
		alu_out = 0;                                    // alu output
		dest_rn = rd;                                   // dest reg number
		wreg    = 0;                                    // write regfile
		wmem    = 0;                                    // write memory (sw)
		rmem    = 0;                                    // read  memory (lw)
		next_pc = pc_plus_4;
		case (1'b1)
			i_add: begin                                // add
				 alu_out = a + b;
				 wreg    = 1; end
			i_addu: begin                               // addu
				 alu_out = a + b;
				 wreg    = 1; end
			i_sub: begin                                // sub
				 alu_out = a - b;
				 wreg    = 1; end
			i_and: begin                                // and
				 alu_out = a & b;
				 wreg    = 1; end
			i_or: begin                                 // or
				 alu_out = a | b;
				 wreg    = 1; end
			i_xor: begin                                // xor
				 alu_out = a ^ b;
				 wreg    = 1; end
			i_sll: begin                                // sll
				 alu_out = b << sa;
				 wreg    = 1; end
			i_srl: begin                                // srl
				 alu_out = b >> sa;
				 wreg    = 1; end
			i_sra: begin                                // sra
				 alu_out = $signed(b) >>> sa;
				 wreg    = 1; end
			i_jr: begin                                 // jr
				 next_pc = a; end
			i_addi: begin                               // addi
				 alu_out = a + {{16{sign}},imm};
				 dest_rn = rt;
				 wreg    = 1; end
			i_addiu: begin                               // addiu
				 alu_out = a + imm;
				 dest_rn = rt;
				 wreg    = 1; end
			i_andi: begin                               // andi
				 alu_out = a & {16'h0,imm};
				 dest_rn = rt;
				 wreg    = 1; end
			i_ori: begin                                // ori
				 alu_out = a | {16'h0,imm};
				 dest_rn = rt;
				 wreg    = 1; end
			i_xori: begin                               // xori
				 alu_out = a ^ {16'h0,imm};
				 dest_rn = rt;
				 wreg    = 1; end
			i_lx:										// lw	// lb	// lbu
				begin                                 
				 alu_out = a + {{16{sign}},imm};
				 dest_rn = rt;
				 rmem    = 1;
				 wreg    = 1; end
			i_sw: begin                                 // sw
				 alu_out = a + {{16{sign}},imm};
				 wmem    = 1; end
			i_beq: begin                                // beq
				 if (a == b) 
					next_pc = pc_plus_4 + offset; end
			i_bne: begin                                // bne
				 if (a != b) 
					next_pc = pc_plus_4 + offset; end
			i_lui: begin                                // lui
				 alu_out = {imm,16'h0};
				 dest_rn = rt;
				 wreg    = 1; end
			i_j: begin                                  // j
				 next_pc = j_addr; end
			i_jal: begin                                // jal
				 alu_out = pc_plus_4;
				 wreg    = 1;
				 dest_rn = 5'd31;
				 next_pc = j_addr; end
			i_slt: begin
				alu_out = $signed(a) < $signed(b) ? 1'b1 : 1'b0;
				wreg = 1;
				dest_rn = rd;
			end
			
			i_slti: begin
				alu_out = $signed(a) < $signed(imm) ? 1'b1 : 1'b0;
				dest_rn = rt;
				wreg	= 1;
			end
			
			
			default: ;
		endcase
	end
endmodule
